-- Lab7.vhd

-- Generated using ACDS version 17.0 595

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Lab7 is
	port (
		clk_clk           : in  std_logic                     := '0';             --        clk.clk
		hex_1_2_export    : out std_logic_vector(13 downto 0);                    --    hex_1_2.export
		hex_3_4_export    : out std_logic_vector(13 downto 0);                    --    hex_3_4.export
		hex_5_6_export    : out std_logic_vector(13 downto 0);                    --    hex_5_6.export
		leds_export       : out std_logic_vector(9 downto 0);                     --       leds.export
		pushbutton_export : in  std_logic_vector(3 downto 0)  := (others => '0'); -- pushbutton.export
		rooms_hex2        : out std_logic_vector(6 downto 0);                     --      rooms.hex2
		rooms_hex1        : out std_logic_vector(6 downto 0);                     --           .hex1
		rooms_hex3        : out std_logic_vector(6 downto 0);                     --           .hex3
		rooms_leds_out    : out std_logic;                                        --           .leds_out
		sw_sliders_export : in  std_logic_vector(9 downto 0)  := (others => '0')  -- sw_sliders.export
	);
end entity Lab7;

architecture rtl of Lab7 is
	component Lab7_Hex_1_2 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(13 downto 0)                     -- export
		);
	end component Lab7_Hex_1_2;

	component Lab7_JTAG_UART is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component Lab7_JTAG_UART;

	component Lab7_MUTEX is
		port (
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			clk           : in  std_logic                     := 'X';             -- clk
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			data_from_cpu : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			read          : in  std_logic                     := 'X';             -- read
			write         : in  std_logic                     := 'X';             -- write
			data_to_cpu   : out std_logic_vector(31 downto 0);                    -- readdata
			address       : in  std_logic                     := 'X'              -- address
		);
	end component Lab7_MUTEX;

	component Lab7_Processor1 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(19 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(19 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component Lab7_Processor1;

	component Lab7_Processor2 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(19 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(19 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component Lab7_Processor2;

	component Lab7_RAM1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component Lab7_RAM1;

	component Lab7_RAM2 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component Lab7_RAM2;

	component Lab7_SHARED_MEMORY is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component Lab7_SHARED_MEMORY;

	component Lab7_Timer1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component Lab7_Timer1;

	component Lab7_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component Lab7_leds;

	component Lab7_pushbutton is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component Lab7_pushbutton;

	component Lab6 is
		port (
			writedata    : in  std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			wr           : in  std_logic                    := 'X';             -- write
			cs           : in  std_logic                    := 'X';             -- chipselect
			hexThree_out : out std_logic_vector(6 downto 0);                    -- hex2
			hexOne_out   : out std_logic_vector(6 downto 0);                    -- hex1
			hexTwo_out   : out std_logic_vector(6 downto 0);                    -- hex3
			leds_out     : out std_logic;                                       -- leds_out
			reset_reset  : in  std_logic                    := 'X';             -- reset
			clk_clk      : in  std_logic                    := 'X'              -- clk
		);
	end component Lab6;

	component Lab7_sw_sliders is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component Lab7_sw_sliders;

	component Lab7_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                    : in  std_logic                     := 'X';             -- clk
			Processor1_reset_reset_bridge_in_reset_reset     : in  std_logic                     := 'X';             -- reset
			Processor2_reset_reset_bridge_in_reset_reset     : in  std_logic                     := 'X';             -- reset
			RAM2_reset1_reset_bridge_in_reset_reset          : in  std_logic                     := 'X';             -- reset
			SHARED_MEMORY_reset1_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			Processor1_data_master_address                   : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			Processor1_data_master_waitrequest               : out std_logic;                                        -- waitrequest
			Processor1_data_master_byteenable                : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			Processor1_data_master_read                      : in  std_logic                     := 'X';             -- read
			Processor1_data_master_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			Processor1_data_master_write                     : in  std_logic                     := 'X';             -- write
			Processor1_data_master_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			Processor1_data_master_debugaccess               : in  std_logic                     := 'X';             -- debugaccess
			Processor1_instruction_master_address            : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			Processor1_instruction_master_waitrequest        : out std_logic;                                        -- waitrequest
			Processor1_instruction_master_read               : in  std_logic                     := 'X';             -- read
			Processor1_instruction_master_readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			Processor2_data_master_address                   : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			Processor2_data_master_waitrequest               : out std_logic;                                        -- waitrequest
			Processor2_data_master_byteenable                : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			Processor2_data_master_read                      : in  std_logic                     := 'X';             -- read
			Processor2_data_master_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			Processor2_data_master_write                     : in  std_logic                     := 'X';             -- write
			Processor2_data_master_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			Processor2_data_master_debugaccess               : in  std_logic                     := 'X';             -- debugaccess
			Processor2_instruction_master_address            : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			Processor2_instruction_master_waitrequest        : out std_logic;                                        -- waitrequest
			Processor2_instruction_master_read               : in  std_logic                     := 'X';             -- read
			Processor2_instruction_master_readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			Hex_1_2_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			Hex_1_2_s1_write                                 : out std_logic;                                        -- write
			Hex_1_2_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Hex_1_2_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			Hex_1_2_s1_chipselect                            : out std_logic;                                        -- chipselect
			Hex_3_4_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			Hex_3_4_s1_write                                 : out std_logic;                                        -- write
			Hex_3_4_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Hex_3_4_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			Hex_3_4_s1_chipselect                            : out std_logic;                                        -- chipselect
			Hex_5_6_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			Hex_5_6_s1_write                                 : out std_logic;                                        -- write
			Hex_5_6_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Hex_5_6_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			Hex_5_6_s1_chipselect                            : out std_logic;                                        -- chipselect
			JTAG_UART_avalon_jtag_slave_address              : out std_logic_vector(0 downto 0);                     -- address
			JTAG_UART_avalon_jtag_slave_write                : out std_logic;                                        -- write
			JTAG_UART_avalon_jtag_slave_read                 : out std_logic;                                        -- read
			JTAG_UART_avalon_jtag_slave_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			JTAG_UART_avalon_jtag_slave_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			JTAG_UART_avalon_jtag_slave_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			JTAG_UART_avalon_jtag_slave_chipselect           : out std_logic;                                        -- chipselect
			leds_s1_address                                  : out std_logic_vector(1 downto 0);                     -- address
			leds_s1_write                                    : out std_logic;                                        -- write
			leds_s1_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			leds_s1_writedata                                : out std_logic_vector(31 downto 0);                    -- writedata
			leds_s1_chipselect                               : out std_logic;                                        -- chipselect
			MUTEX_s1_address                                 : out std_logic_vector(0 downto 0);                     -- address
			MUTEX_s1_write                                   : out std_logic;                                        -- write
			MUTEX_s1_read                                    : out std_logic;                                        -- read
			MUTEX_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			MUTEX_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			MUTEX_s1_chipselect                              : out std_logic;                                        -- chipselect
			Processor1_debug_mem_slave_address               : out std_logic_vector(8 downto 0);                     -- address
			Processor1_debug_mem_slave_write                 : out std_logic;                                        -- write
			Processor1_debug_mem_slave_read                  : out std_logic;                                        -- read
			Processor1_debug_mem_slave_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Processor1_debug_mem_slave_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			Processor1_debug_mem_slave_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			Processor1_debug_mem_slave_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			Processor1_debug_mem_slave_debugaccess           : out std_logic;                                        -- debugaccess
			Processor2_debug_mem_slave_address               : out std_logic_vector(8 downto 0);                     -- address
			Processor2_debug_mem_slave_write                 : out std_logic;                                        -- write
			Processor2_debug_mem_slave_read                  : out std_logic;                                        -- read
			Processor2_debug_mem_slave_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Processor2_debug_mem_slave_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			Processor2_debug_mem_slave_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			Processor2_debug_mem_slave_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			Processor2_debug_mem_slave_debugaccess           : out std_logic;                                        -- debugaccess
			pushbutton_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			pushbutton_s1_write                              : out std_logic;                                        -- write
			pushbutton_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pushbutton_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			pushbutton_s1_chipselect                         : out std_logic;                                        -- chipselect
			RAM1_s1_address                                  : out std_logic_vector(15 downto 0);                    -- address
			RAM1_s1_write                                    : out std_logic;                                        -- write
			RAM1_s1_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			RAM1_s1_writedata                                : out std_logic_vector(31 downto 0);                    -- writedata
			RAM1_s1_byteenable                               : out std_logic_vector(3 downto 0);                     -- byteenable
			RAM1_s1_chipselect                               : out std_logic;                                        -- chipselect
			RAM1_s1_clken                                    : out std_logic;                                        -- clken
			RAM2_s1_address                                  : out std_logic_vector(14 downto 0);                    -- address
			RAM2_s1_write                                    : out std_logic;                                        -- write
			RAM2_s1_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			RAM2_s1_writedata                                : out std_logic_vector(31 downto 0);                    -- writedata
			RAM2_s1_byteenable                               : out std_logic_vector(3 downto 0);                     -- byteenable
			RAM2_s1_chipselect                               : out std_logic;                                        -- chipselect
			RAM2_s1_clken                                    : out std_logic;                                        -- clken
			rooms_manager_0_avalon_slave_0_write             : out std_logic;                                        -- write
			rooms_manager_0_avalon_slave_0_writedata         : out std_logic_vector(7 downto 0);                     -- writedata
			rooms_manager_0_avalon_slave_0_chipselect        : out std_logic;                                        -- chipselect
			SHARED_MEMORY_s1_address                         : out std_logic_vector(9 downto 0);                     -- address
			SHARED_MEMORY_s1_write                           : out std_logic;                                        -- write
			SHARED_MEMORY_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			SHARED_MEMORY_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			SHARED_MEMORY_s1_byteenable                      : out std_logic_vector(3 downto 0);                     -- byteenable
			SHARED_MEMORY_s1_chipselect                      : out std_logic;                                        -- chipselect
			SHARED_MEMORY_s1_clken                           : out std_logic;                                        -- clken
			sw_sliders_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			sw_sliders_s1_write                              : out std_logic;                                        -- write
			sw_sliders_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sw_sliders_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			sw_sliders_s1_chipselect                         : out std_logic;                                        -- chipselect
			Timer1_s1_address                                : out std_logic_vector(2 downto 0);                     -- address
			Timer1_s1_write                                  : out std_logic;                                        -- write
			Timer1_s1_readdata                               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			Timer1_s1_writedata                              : out std_logic_vector(15 downto 0);                    -- writedata
			Timer1_s1_chipselect                             : out std_logic;                                        -- chipselect
			Timer2_s1_address                                : out std_logic_vector(2 downto 0);                     -- address
			Timer2_s1_write                                  : out std_logic;                                        -- write
			Timer2_s1_readdata                               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			Timer2_s1_writedata                              : out std_logic_vector(15 downto 0);                    -- writedata
			Timer2_s1_chipselect                             : out std_logic                                         -- chipselect
		);
	end component Lab7_mm_interconnect_0;

	component Lab7_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component Lab7_irq_mapper;

	component Lab7_irq_mapper_001 is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component Lab7_irq_mapper_001;

	component lab7_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component lab7_rst_controller;

	component lab7_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			reset_in2      : in  std_logic := 'X'; -- reset_in2.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component lab7_rst_controller_001;

	component lab7_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component lab7_rst_controller_002;

	signal processor1_debug_reset_request_reset                          : std_logic;                     -- Processor1:debug_reset_request -> [rst_controller:reset_in0, rst_controller:reset_in1, rst_controller_001:reset_in0, rst_controller_001:reset_in2, rst_controller_002:reset_in0, rst_controller_003:reset_in0]
	signal processor1_data_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:Processor1_data_master_readdata -> Processor1:d_readdata
	signal processor1_data_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:Processor1_data_master_waitrequest -> Processor1:d_waitrequest
	signal processor1_data_master_debugaccess                            : std_logic;                     -- Processor1:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Processor1_data_master_debugaccess
	signal processor1_data_master_address                                : std_logic_vector(19 downto 0); -- Processor1:d_address -> mm_interconnect_0:Processor1_data_master_address
	signal processor1_data_master_byteenable                             : std_logic_vector(3 downto 0);  -- Processor1:d_byteenable -> mm_interconnect_0:Processor1_data_master_byteenable
	signal processor1_data_master_read                                   : std_logic;                     -- Processor1:d_read -> mm_interconnect_0:Processor1_data_master_read
	signal processor1_data_master_write                                  : std_logic;                     -- Processor1:d_write -> mm_interconnect_0:Processor1_data_master_write
	signal processor1_data_master_writedata                              : std_logic_vector(31 downto 0); -- Processor1:d_writedata -> mm_interconnect_0:Processor1_data_master_writedata
	signal processor2_data_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:Processor2_data_master_readdata -> Processor2:d_readdata
	signal processor2_data_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:Processor2_data_master_waitrequest -> Processor2:d_waitrequest
	signal processor2_data_master_debugaccess                            : std_logic;                     -- Processor2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Processor2_data_master_debugaccess
	signal processor2_data_master_address                                : std_logic_vector(19 downto 0); -- Processor2:d_address -> mm_interconnect_0:Processor2_data_master_address
	signal processor2_data_master_byteenable                             : std_logic_vector(3 downto 0);  -- Processor2:d_byteenable -> mm_interconnect_0:Processor2_data_master_byteenable
	signal processor2_data_master_read                                   : std_logic;                     -- Processor2:d_read -> mm_interconnect_0:Processor2_data_master_read
	signal processor2_data_master_write                                  : std_logic;                     -- Processor2:d_write -> mm_interconnect_0:Processor2_data_master_write
	signal processor2_data_master_writedata                              : std_logic_vector(31 downto 0); -- Processor2:d_writedata -> mm_interconnect_0:Processor2_data_master_writedata
	signal processor2_instruction_master_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:Processor2_instruction_master_readdata -> Processor2:i_readdata
	signal processor2_instruction_master_waitrequest                     : std_logic;                     -- mm_interconnect_0:Processor2_instruction_master_waitrequest -> Processor2:i_waitrequest
	signal processor2_instruction_master_address                         : std_logic_vector(19 downto 0); -- Processor2:i_address -> mm_interconnect_0:Processor2_instruction_master_address
	signal processor2_instruction_master_read                            : std_logic;                     -- Processor2:i_read -> mm_interconnect_0:Processor2_instruction_master_read
	signal processor1_instruction_master_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:Processor1_instruction_master_readdata -> Processor1:i_readdata
	signal processor1_instruction_master_waitrequest                     : std_logic;                     -- mm_interconnect_0:Processor1_instruction_master_waitrequest -> Processor1:i_waitrequest
	signal processor1_instruction_master_address                         : std_logic_vector(19 downto 0); -- Processor1:i_address -> mm_interconnect_0:Processor1_instruction_master_address
	signal processor1_instruction_master_read                            : std_logic;                     -- Processor1:i_read -> mm_interconnect_0:Processor1_instruction_master_read
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	signal mm_interconnect_0_processor1_debug_mem_slave_readdata         : std_logic_vector(31 downto 0); -- Processor1:debug_mem_slave_readdata -> mm_interconnect_0:Processor1_debug_mem_slave_readdata
	signal mm_interconnect_0_processor1_debug_mem_slave_waitrequest      : std_logic;                     -- Processor1:debug_mem_slave_waitrequest -> mm_interconnect_0:Processor1_debug_mem_slave_waitrequest
	signal mm_interconnect_0_processor1_debug_mem_slave_debugaccess      : std_logic;                     -- mm_interconnect_0:Processor1_debug_mem_slave_debugaccess -> Processor1:debug_mem_slave_debugaccess
	signal mm_interconnect_0_processor1_debug_mem_slave_address          : std_logic_vector(8 downto 0);  -- mm_interconnect_0:Processor1_debug_mem_slave_address -> Processor1:debug_mem_slave_address
	signal mm_interconnect_0_processor1_debug_mem_slave_read             : std_logic;                     -- mm_interconnect_0:Processor1_debug_mem_slave_read -> Processor1:debug_mem_slave_read
	signal mm_interconnect_0_processor1_debug_mem_slave_byteenable       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Processor1_debug_mem_slave_byteenable -> Processor1:debug_mem_slave_byteenable
	signal mm_interconnect_0_processor1_debug_mem_slave_write            : std_logic;                     -- mm_interconnect_0:Processor1_debug_mem_slave_write -> Processor1:debug_mem_slave_write
	signal mm_interconnect_0_processor1_debug_mem_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:Processor1_debug_mem_slave_writedata -> Processor1:debug_mem_slave_writedata
	signal mm_interconnect_0_ram1_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:RAM1_s1_chipselect -> RAM1:chipselect
	signal mm_interconnect_0_ram1_s1_readdata                            : std_logic_vector(31 downto 0); -- RAM1:readdata -> mm_interconnect_0:RAM1_s1_readdata
	signal mm_interconnect_0_ram1_s1_address                             : std_logic_vector(15 downto 0); -- mm_interconnect_0:RAM1_s1_address -> RAM1:address
	signal mm_interconnect_0_ram1_s1_byteenable                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:RAM1_s1_byteenable -> RAM1:byteenable
	signal mm_interconnect_0_ram1_s1_write                               : std_logic;                     -- mm_interconnect_0:RAM1_s1_write -> RAM1:write
	signal mm_interconnect_0_ram1_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:RAM1_s1_writedata -> RAM1:writedata
	signal mm_interconnect_0_ram1_s1_clken                               : std_logic;                     -- mm_interconnect_0:RAM1_s1_clken -> RAM1:clken
	signal mm_interconnect_0_sw_sliders_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:sw_sliders_s1_chipselect -> sw_sliders:chipselect
	signal mm_interconnect_0_sw_sliders_s1_readdata                      : std_logic_vector(31 downto 0); -- sw_sliders:readdata -> mm_interconnect_0:sw_sliders_s1_readdata
	signal mm_interconnect_0_sw_sliders_s1_address                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sw_sliders_s1_address -> sw_sliders:address
	signal mm_interconnect_0_sw_sliders_s1_write                         : std_logic;                     -- mm_interconnect_0:sw_sliders_s1_write -> mm_interconnect_0_sw_sliders_s1_write:in
	signal mm_interconnect_0_sw_sliders_s1_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:sw_sliders_s1_writedata -> sw_sliders:writedata
	signal mm_interconnect_0_timer1_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:Timer1_s1_chipselect -> Timer1:chipselect
	signal mm_interconnect_0_timer1_s1_readdata                          : std_logic_vector(15 downto 0); -- Timer1:readdata -> mm_interconnect_0:Timer1_s1_readdata
	signal mm_interconnect_0_timer1_s1_address                           : std_logic_vector(2 downto 0);  -- mm_interconnect_0:Timer1_s1_address -> Timer1:address
	signal mm_interconnect_0_timer1_s1_write                             : std_logic;                     -- mm_interconnect_0:Timer1_s1_write -> mm_interconnect_0_timer1_s1_write:in
	signal mm_interconnect_0_timer1_s1_writedata                         : std_logic_vector(15 downto 0); -- mm_interconnect_0:Timer1_s1_writedata -> Timer1:writedata
	signal mm_interconnect_0_shared_memory_s1_chipselect                 : std_logic;                     -- mm_interconnect_0:SHARED_MEMORY_s1_chipselect -> SHARED_MEMORY:chipselect
	signal mm_interconnect_0_shared_memory_s1_readdata                   : std_logic_vector(31 downto 0); -- SHARED_MEMORY:readdata -> mm_interconnect_0:SHARED_MEMORY_s1_readdata
	signal mm_interconnect_0_shared_memory_s1_address                    : std_logic_vector(9 downto 0);  -- mm_interconnect_0:SHARED_MEMORY_s1_address -> SHARED_MEMORY:address
	signal mm_interconnect_0_shared_memory_s1_byteenable                 : std_logic_vector(3 downto 0);  -- mm_interconnect_0:SHARED_MEMORY_s1_byteenable -> SHARED_MEMORY:byteenable
	signal mm_interconnect_0_shared_memory_s1_write                      : std_logic;                     -- mm_interconnect_0:SHARED_MEMORY_s1_write -> SHARED_MEMORY:write
	signal mm_interconnect_0_shared_memory_s1_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:SHARED_MEMORY_s1_writedata -> SHARED_MEMORY:writedata
	signal mm_interconnect_0_shared_memory_s1_clken                      : std_logic;                     -- mm_interconnect_0:SHARED_MEMORY_s1_clken -> SHARED_MEMORY:clken
	signal mm_interconnect_0_mutex_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:MUTEX_s1_chipselect -> MUTEX:chipselect
	signal mm_interconnect_0_mutex_s1_readdata                           : std_logic_vector(31 downto 0); -- MUTEX:data_to_cpu -> mm_interconnect_0:MUTEX_s1_readdata
	signal mm_interconnect_0_mutex_s1_address                            : std_logic_vector(0 downto 0);  -- mm_interconnect_0:MUTEX_s1_address -> MUTEX:address
	signal mm_interconnect_0_mutex_s1_read                               : std_logic;                     -- mm_interconnect_0:MUTEX_s1_read -> MUTEX:read
	signal mm_interconnect_0_mutex_s1_write                              : std_logic;                     -- mm_interconnect_0:MUTEX_s1_write -> MUTEX:write
	signal mm_interconnect_0_mutex_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:MUTEX_s1_writedata -> MUTEX:data_from_cpu
	signal mm_interconnect_0_pushbutton_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:pushbutton_s1_chipselect -> pushbutton:chipselect
	signal mm_interconnect_0_pushbutton_s1_readdata                      : std_logic_vector(31 downto 0); -- pushbutton:readdata -> mm_interconnect_0:pushbutton_s1_readdata
	signal mm_interconnect_0_pushbutton_s1_address                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pushbutton_s1_address -> pushbutton:address
	signal mm_interconnect_0_pushbutton_s1_write                         : std_logic;                     -- mm_interconnect_0:pushbutton_s1_write -> mm_interconnect_0_pushbutton_s1_write:in
	signal mm_interconnect_0_pushbutton_s1_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:pushbutton_s1_writedata -> pushbutton:writedata
	signal mm_interconnect_0_processor2_debug_mem_slave_readdata         : std_logic_vector(31 downto 0); -- Processor2:debug_mem_slave_readdata -> mm_interconnect_0:Processor2_debug_mem_slave_readdata
	signal mm_interconnect_0_processor2_debug_mem_slave_waitrequest      : std_logic;                     -- Processor2:debug_mem_slave_waitrequest -> mm_interconnect_0:Processor2_debug_mem_slave_waitrequest
	signal mm_interconnect_0_processor2_debug_mem_slave_debugaccess      : std_logic;                     -- mm_interconnect_0:Processor2_debug_mem_slave_debugaccess -> Processor2:debug_mem_slave_debugaccess
	signal mm_interconnect_0_processor2_debug_mem_slave_address          : std_logic_vector(8 downto 0);  -- mm_interconnect_0:Processor2_debug_mem_slave_address -> Processor2:debug_mem_slave_address
	signal mm_interconnect_0_processor2_debug_mem_slave_read             : std_logic;                     -- mm_interconnect_0:Processor2_debug_mem_slave_read -> Processor2:debug_mem_slave_read
	signal mm_interconnect_0_processor2_debug_mem_slave_byteenable       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Processor2_debug_mem_slave_byteenable -> Processor2:debug_mem_slave_byteenable
	signal mm_interconnect_0_processor2_debug_mem_slave_write            : std_logic;                     -- mm_interconnect_0:Processor2_debug_mem_slave_write -> Processor2:debug_mem_slave_write
	signal mm_interconnect_0_processor2_debug_mem_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:Processor2_debug_mem_slave_writedata -> Processor2:debug_mem_slave_writedata
	signal mm_interconnect_0_ram2_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:RAM2_s1_chipselect -> RAM2:chipselect
	signal mm_interconnect_0_ram2_s1_readdata                            : std_logic_vector(31 downto 0); -- RAM2:readdata -> mm_interconnect_0:RAM2_s1_readdata
	signal mm_interconnect_0_ram2_s1_address                             : std_logic_vector(14 downto 0); -- mm_interconnect_0:RAM2_s1_address -> RAM2:address
	signal mm_interconnect_0_ram2_s1_byteenable                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:RAM2_s1_byteenable -> RAM2:byteenable
	signal mm_interconnect_0_ram2_s1_write                               : std_logic;                     -- mm_interconnect_0:RAM2_s1_write -> RAM2:write
	signal mm_interconnect_0_ram2_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:RAM2_s1_writedata -> RAM2:writedata
	signal mm_interconnect_0_ram2_s1_clken                               : std_logic;                     -- mm_interconnect_0:RAM2_s1_clken -> RAM2:clken
	signal mm_interconnect_0_timer2_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:Timer2_s1_chipselect -> Timer2:chipselect
	signal mm_interconnect_0_timer2_s1_readdata                          : std_logic_vector(15 downto 0); -- Timer2:readdata -> mm_interconnect_0:Timer2_s1_readdata
	signal mm_interconnect_0_timer2_s1_address                           : std_logic_vector(2 downto 0);  -- mm_interconnect_0:Timer2_s1_address -> Timer2:address
	signal mm_interconnect_0_timer2_s1_write                             : std_logic;                     -- mm_interconnect_0:Timer2_s1_write -> mm_interconnect_0_timer2_s1_write:in
	signal mm_interconnect_0_timer2_s1_writedata                         : std_logic_vector(15 downto 0); -- mm_interconnect_0:Timer2_s1_writedata -> Timer2:writedata
	signal mm_interconnect_0_hex_5_6_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:Hex_5_6_s1_chipselect -> Hex_5_6:chipselect
	signal mm_interconnect_0_hex_5_6_s1_readdata                         : std_logic_vector(31 downto 0); -- Hex_5_6:readdata -> mm_interconnect_0:Hex_5_6_s1_readdata
	signal mm_interconnect_0_hex_5_6_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Hex_5_6_s1_address -> Hex_5_6:address
	signal mm_interconnect_0_hex_5_6_s1_write                            : std_logic;                     -- mm_interconnect_0:Hex_5_6_s1_write -> mm_interconnect_0_hex_5_6_s1_write:in
	signal mm_interconnect_0_hex_5_6_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:Hex_5_6_s1_writedata -> Hex_5_6:writedata
	signal mm_interconnect_0_hex_3_4_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:Hex_3_4_s1_chipselect -> Hex_3_4:chipselect
	signal mm_interconnect_0_hex_3_4_s1_readdata                         : std_logic_vector(31 downto 0); -- Hex_3_4:readdata -> mm_interconnect_0:Hex_3_4_s1_readdata
	signal mm_interconnect_0_hex_3_4_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Hex_3_4_s1_address -> Hex_3_4:address
	signal mm_interconnect_0_hex_3_4_s1_write                            : std_logic;                     -- mm_interconnect_0:Hex_3_4_s1_write -> mm_interconnect_0_hex_3_4_s1_write:in
	signal mm_interconnect_0_hex_3_4_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:Hex_3_4_s1_writedata -> Hex_3_4:writedata
	signal mm_interconnect_0_hex_1_2_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:Hex_1_2_s1_chipselect -> Hex_1_2:chipselect
	signal mm_interconnect_0_hex_1_2_s1_readdata                         : std_logic_vector(31 downto 0); -- Hex_1_2:readdata -> mm_interconnect_0:Hex_1_2_s1_readdata
	signal mm_interconnect_0_hex_1_2_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Hex_1_2_s1_address -> Hex_1_2:address
	signal mm_interconnect_0_hex_1_2_s1_write                            : std_logic;                     -- mm_interconnect_0:Hex_1_2_s1_write -> mm_interconnect_0_hex_1_2_s1_write:in
	signal mm_interconnect_0_hex_1_2_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:Hex_1_2_s1_writedata -> Hex_1_2:writedata
	signal mm_interconnect_0_leds_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	signal mm_interconnect_0_leds_s1_readdata                            : std_logic_vector(31 downto 0); -- leds:readdata -> mm_interconnect_0:leds_s1_readdata
	signal mm_interconnect_0_leds_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:leds_s1_address -> leds:address
	signal mm_interconnect_0_leds_s1_write                               : std_logic;                     -- mm_interconnect_0:leds_s1_write -> mm_interconnect_0_leds_s1_write:in
	signal mm_interconnect_0_leds_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:leds_s1_writedata -> leds:writedata
	signal mm_interconnect_0_rooms_manager_0_avalon_slave_0_chipselect   : std_logic;                     -- mm_interconnect_0:rooms_manager_0_avalon_slave_0_chipselect -> rooms_manager_0:cs
	signal mm_interconnect_0_rooms_manager_0_avalon_slave_0_write        : std_logic;                     -- mm_interconnect_0:rooms_manager_0_avalon_slave_0_write -> rooms_manager_0:wr
	signal mm_interconnect_0_rooms_manager_0_avalon_slave_0_writedata    : std_logic_vector(7 downto 0);  -- mm_interconnect_0:rooms_manager_0_avalon_slave_0_writedata -> rooms_manager_0:writedata
	signal irq_mapper_receiver3_irq                                      : std_logic;                     -- Timer1:irq -> irq_mapper:receiver3_irq
	signal processor1_irq_irq                                            : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> Processor1:irq
	signal irq_mapper_001_receiver0_irq                                  : std_logic;                     -- Timer2:irq -> irq_mapper_001:receiver0_irq
	signal processor2_irq_irq                                            : std_logic_vector(31 downto 0); -- irq_mapper_001:sender_irq -> Processor2:irq
	signal irq_mapper_receiver2_irq                                      : std_logic;                     -- JTAG_UART:av_irq -> [irq_mapper:receiver2_irq, irq_mapper_001:receiver3_irq]
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- pushbutton:irq -> [irq_mapper:receiver1_irq, irq_mapper_001:receiver1_irq]
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- sw_sliders:irq -> [irq_mapper:receiver0_irq, irq_mapper_001:receiver2_irq]
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [RAM1:reset, irq_mapper:reset, mm_interconnect_0:Processor1_reset_reset_bridge_in_reset_reset, rooms_manager_0:reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                            : std_logic;                     -- rst_controller:reset_req -> [Processor1:reset_req, RAM1:reset_req, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                            : std_logic;                     -- rst_controller_001:reset_out -> [SHARED_MEMORY:reset, mm_interconnect_0:SHARED_MEMORY_reset1_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset_req                        : std_logic;                     -- rst_controller_001:reset_req -> [SHARED_MEMORY:reset_req, rst_translator_001:reset_req_in]
	signal processor2_debug_reset_request_reset                          : std_logic;                     -- Processor2:debug_reset_request -> [rst_controller_001:reset_in1, rst_controller_003:reset_in1]
	signal rst_controller_002_reset_out_reset                            : std_logic;                     -- rst_controller_002:reset_out -> [irq_mapper_001:reset, mm_interconnect_0:Processor2_reset_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in]
	signal rst_controller_002_reset_out_reset_req                        : std_logic;                     -- rst_controller_002:reset_req -> [Processor2:reset_req, rst_translator_002:reset_req_in]
	signal rst_controller_003_reset_out_reset                            : std_logic;                     -- rst_controller_003:reset_out -> [RAM2:reset, mm_interconnect_0:RAM2_reset1_reset_bridge_in_reset_reset, rst_controller_003_reset_out_reset:in]
	signal rst_controller_003_reset_out_reset_req                        : std_logic;                     -- rst_controller_003:reset_req -> [RAM2:reset_req, rst_translator_003:reset_req_in]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> JTAG_UART:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> JTAG_UART:av_write_n
	signal mm_interconnect_0_sw_sliders_s1_write_ports_inv               : std_logic;                     -- mm_interconnect_0_sw_sliders_s1_write:inv -> sw_sliders:write_n
	signal mm_interconnect_0_timer1_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_timer1_s1_write:inv -> Timer1:write_n
	signal mm_interconnect_0_pushbutton_s1_write_ports_inv               : std_logic;                     -- mm_interconnect_0_pushbutton_s1_write:inv -> pushbutton:write_n
	signal mm_interconnect_0_timer2_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_timer2_s1_write:inv -> Timer2:write_n
	signal mm_interconnect_0_hex_5_6_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_hex_5_6_s1_write:inv -> Hex_5_6:write_n
	signal mm_interconnect_0_hex_3_4_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_hex_3_4_s1_write:inv -> Hex_3_4:write_n
	signal mm_interconnect_0_hex_1_2_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_hex_1_2_s1_write:inv -> Hex_1_2:write_n
	signal mm_interconnect_0_leds_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_leds_s1_write:inv -> leds:write_n
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [Hex_1_2:reset_n, Hex_3_4:reset_n, Hex_5_6:reset_n, JTAG_UART:rst_n, Processor1:reset_n, Timer1:reset_n, leds:reset_n, pushbutton:reset_n, sw_sliders:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> MUTEX:reset_n
	signal rst_controller_002_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> Processor2:reset_n
	signal rst_controller_003_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_003_reset_out_reset:inv -> Timer2:reset_n

begin

	hex_1_2 : component Lab7_Hex_1_2
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_hex_1_2_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_1_2_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_1_2_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_1_2_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_1_2_s1_readdata,        --                    .readdata
			out_port   => hex_1_2_export                                -- external_connection.export
		);

	hex_3_4 : component Lab7_Hex_1_2
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_hex_3_4_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_3_4_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_3_4_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_3_4_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_3_4_s1_readdata,        --                    .readdata
			out_port   => hex_3_4_export                                -- external_connection.export
		);

	hex_5_6 : component Lab7_Hex_1_2
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_hex_5_6_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_5_6_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_5_6_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_5_6_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_5_6_s1_readdata,        --                    .readdata
			out_port   => hex_5_6_export                                -- external_connection.export
		);

	jtag_uart : component Lab7_JTAG_UART
		port map (
			clk            => clk_clk,                                                       --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver2_irq                                       --               irq.irq
		);

	mutex : component Lab7_MUTEX
		port map (
			reset_n       => rst_controller_001_reset_out_reset_ports_inv, -- reset.reset_n
			clk           => clk_clk,                                      --   clk.clk
			chipselect    => mm_interconnect_0_mutex_s1_chipselect,        --    s1.chipselect
			data_from_cpu => mm_interconnect_0_mutex_s1_writedata,         --      .writedata
			read          => mm_interconnect_0_mutex_s1_read,              --      .read
			write         => mm_interconnect_0_mutex_s1_write,             --      .write
			data_to_cpu   => mm_interconnect_0_mutex_s1_readdata,          --      .readdata
			address       => mm_interconnect_0_mutex_s1_address(0)         --      .address
		);

	processor1 : component Lab7_Processor1
		port map (
			clk                                 => clk_clk,                                                  --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                 --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                       --                          .reset_req
			d_address                           => processor1_data_master_address,                           --               data_master.address
			d_byteenable                        => processor1_data_master_byteenable,                        --                          .byteenable
			d_read                              => processor1_data_master_read,                              --                          .read
			d_readdata                          => processor1_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => processor1_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => processor1_data_master_write,                             --                          .write
			d_writedata                         => processor1_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => processor1_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => processor1_instruction_master_address,                    --        instruction_master.address
			i_read                              => processor1_instruction_master_read,                       --                          .read
			i_readdata                          => processor1_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => processor1_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => processor1_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => processor1_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_processor1_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_processor1_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_processor1_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_processor1_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_processor1_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_processor1_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_processor1_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_processor1_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                      -- custom_instruction_master.readra
		);

	processor2 : component Lab7_Processor2
		port map (
			clk                                 => clk_clk,                                                  --                       clk.clk
			reset_n                             => rst_controller_002_reset_out_reset_ports_inv,             --                     reset.reset_n
			reset_req                           => rst_controller_002_reset_out_reset_req,                   --                          .reset_req
			d_address                           => processor2_data_master_address,                           --               data_master.address
			d_byteenable                        => processor2_data_master_byteenable,                        --                          .byteenable
			d_read                              => processor2_data_master_read,                              --                          .read
			d_readdata                          => processor2_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => processor2_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => processor2_data_master_write,                             --                          .write
			d_writedata                         => processor2_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => processor2_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => processor2_instruction_master_address,                    --        instruction_master.address
			i_read                              => processor2_instruction_master_read,                       --                          .read
			i_readdata                          => processor2_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => processor2_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => processor2_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => processor2_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_processor2_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_processor2_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_processor2_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_processor2_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_processor2_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_processor2_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_processor2_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_processor2_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                      -- custom_instruction_master.readra
		);

	ram1 : component Lab7_RAM1
		port map (
			clk        => clk_clk,                              --   clk1.clk
			address    => mm_interconnect_0_ram1_s1_address,    --     s1.address
			clken      => mm_interconnect_0_ram1_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_ram1_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_ram1_s1_write,      --       .write
			readdata   => mm_interconnect_0_ram1_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_ram1_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_ram1_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,       -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,   --       .reset_req
			freeze     => '0'                                   -- (terminated)
		);

	ram2 : component Lab7_RAM2
		port map (
			clk        => clk_clk,                                --   clk1.clk
			address    => mm_interconnect_0_ram2_s1_address,      --     s1.address
			clken      => mm_interconnect_0_ram2_s1_clken,        --       .clken
			chipselect => mm_interconnect_0_ram2_s1_chipselect,   --       .chipselect
			write      => mm_interconnect_0_ram2_s1_write,        --       .write
			readdata   => mm_interconnect_0_ram2_s1_readdata,     --       .readdata
			writedata  => mm_interconnect_0_ram2_s1_writedata,    --       .writedata
			byteenable => mm_interconnect_0_ram2_s1_byteenable,   --       .byteenable
			reset      => rst_controller_003_reset_out_reset,     -- reset1.reset
			reset_req  => rst_controller_003_reset_out_reset_req, --       .reset_req
			freeze     => '0'                                     -- (terminated)
		);

	shared_memory : component Lab7_SHARED_MEMORY
		port map (
			clk        => clk_clk,                                       --   clk1.clk
			address    => mm_interconnect_0_shared_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_0_shared_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_shared_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_shared_memory_s1_write,      --       .write
			readdata   => mm_interconnect_0_shared_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_shared_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_shared_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_001_reset_out_reset,            -- reset1.reset
			reset_req  => rst_controller_001_reset_out_reset_req,        --       .reset_req
			freeze     => '0'                                            -- (terminated)
		);

	timer1 : component Lab7_Timer1
		port map (
			clk        => clk_clk,                                     --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    -- reset.reset_n
			address    => mm_interconnect_0_timer1_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer1_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer1_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer1_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer1_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver3_irq                     --   irq.irq
		);

	timer2 : component Lab7_Timer1
		port map (
			clk        => clk_clk,                                      --   clk.clk
			reset_n    => rst_controller_003_reset_out_reset_ports_inv, -- reset.reset_n
			address    => mm_interconnect_0_timer2_s1_address,          --    s1.address
			writedata  => mm_interconnect_0_timer2_s1_writedata,        --      .writedata
			readdata   => mm_interconnect_0_timer2_s1_readdata,         --      .readdata
			chipselect => mm_interconnect_0_timer2_s1_chipselect,       --      .chipselect
			write_n    => mm_interconnect_0_timer2_s1_write_ports_inv,  --      .write_n
			irq        => irq_mapper_001_receiver0_irq                  --   irq.irq
		);

	leds : component Lab7_leds
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_leds_s1_readdata,        --                    .readdata
			out_port   => leds_export                                -- external_connection.export
		);

	pushbutton : component Lab7_pushbutton
		port map (
			clk        => clk_clk,                                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_0_pushbutton_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pushbutton_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pushbutton_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pushbutton_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pushbutton_s1_readdata,        --                    .readdata
			in_port    => pushbutton_export,                               -- external_connection.export
			irq        => irq_mapper_receiver1_irq                         --                 irq.irq
		);

	rooms_manager_0 : component Lab6
		port map (
			writedata    => mm_interconnect_0_rooms_manager_0_avalon_slave_0_writedata,  -- avalon_slave_0.writedata
			wr           => mm_interconnect_0_rooms_manager_0_avalon_slave_0_write,      --               .write
			cs           => mm_interconnect_0_rooms_manager_0_avalon_slave_0_chipselect, --               .chipselect
			hexThree_out => rooms_hex2,                                                  --    conduit_end.hex2
			hexOne_out   => rooms_hex1,                                                  --               .hex1
			hexTwo_out   => rooms_hex3,                                                  --               .hex3
			leds_out     => rooms_leds_out,                                              --               .leds_out
			reset_reset  => rst_controller_reset_out_reset,                              --    reset_reset.reset
			clk_clk      => clk_clk                                                      --        clk_clk.clk
		);

	sw_sliders : component Lab7_sw_sliders
		port map (
			clk        => clk_clk,                                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_0_sw_sliders_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_sw_sliders_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_sw_sliders_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_sw_sliders_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_sw_sliders_s1_readdata,        --                    .readdata
			in_port    => sw_sliders_export,                               -- external_connection.export
			irq        => irq_mapper_receiver0_irq                         --                 irq.irq
		);

	mm_interconnect_0 : component Lab7_mm_interconnect_0
		port map (
			clk_0_clk_clk                                    => clk_clk,                                                     --                                  clk_0_clk.clk
			Processor1_reset_reset_bridge_in_reset_reset     => rst_controller_reset_out_reset,                              --     Processor1_reset_reset_bridge_in_reset.reset
			Processor2_reset_reset_bridge_in_reset_reset     => rst_controller_002_reset_out_reset,                          --     Processor2_reset_reset_bridge_in_reset.reset
			RAM2_reset1_reset_bridge_in_reset_reset          => rst_controller_003_reset_out_reset,                          --          RAM2_reset1_reset_bridge_in_reset.reset
			SHARED_MEMORY_reset1_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                          -- SHARED_MEMORY_reset1_reset_bridge_in_reset.reset
			Processor1_data_master_address                   => processor1_data_master_address,                              --                     Processor1_data_master.address
			Processor1_data_master_waitrequest               => processor1_data_master_waitrequest,                          --                                           .waitrequest
			Processor1_data_master_byteenable                => processor1_data_master_byteenable,                           --                                           .byteenable
			Processor1_data_master_read                      => processor1_data_master_read,                                 --                                           .read
			Processor1_data_master_readdata                  => processor1_data_master_readdata,                             --                                           .readdata
			Processor1_data_master_write                     => processor1_data_master_write,                                --                                           .write
			Processor1_data_master_writedata                 => processor1_data_master_writedata,                            --                                           .writedata
			Processor1_data_master_debugaccess               => processor1_data_master_debugaccess,                          --                                           .debugaccess
			Processor1_instruction_master_address            => processor1_instruction_master_address,                       --              Processor1_instruction_master.address
			Processor1_instruction_master_waitrequest        => processor1_instruction_master_waitrequest,                   --                                           .waitrequest
			Processor1_instruction_master_read               => processor1_instruction_master_read,                          --                                           .read
			Processor1_instruction_master_readdata           => processor1_instruction_master_readdata,                      --                                           .readdata
			Processor2_data_master_address                   => processor2_data_master_address,                              --                     Processor2_data_master.address
			Processor2_data_master_waitrequest               => processor2_data_master_waitrequest,                          --                                           .waitrequest
			Processor2_data_master_byteenable                => processor2_data_master_byteenable,                           --                                           .byteenable
			Processor2_data_master_read                      => processor2_data_master_read,                                 --                                           .read
			Processor2_data_master_readdata                  => processor2_data_master_readdata,                             --                                           .readdata
			Processor2_data_master_write                     => processor2_data_master_write,                                --                                           .write
			Processor2_data_master_writedata                 => processor2_data_master_writedata,                            --                                           .writedata
			Processor2_data_master_debugaccess               => processor2_data_master_debugaccess,                          --                                           .debugaccess
			Processor2_instruction_master_address            => processor2_instruction_master_address,                       --              Processor2_instruction_master.address
			Processor2_instruction_master_waitrequest        => processor2_instruction_master_waitrequest,                   --                                           .waitrequest
			Processor2_instruction_master_read               => processor2_instruction_master_read,                          --                                           .read
			Processor2_instruction_master_readdata           => processor2_instruction_master_readdata,                      --                                           .readdata
			Hex_1_2_s1_address                               => mm_interconnect_0_hex_1_2_s1_address,                        --                                 Hex_1_2_s1.address
			Hex_1_2_s1_write                                 => mm_interconnect_0_hex_1_2_s1_write,                          --                                           .write
			Hex_1_2_s1_readdata                              => mm_interconnect_0_hex_1_2_s1_readdata,                       --                                           .readdata
			Hex_1_2_s1_writedata                             => mm_interconnect_0_hex_1_2_s1_writedata,                      --                                           .writedata
			Hex_1_2_s1_chipselect                            => mm_interconnect_0_hex_1_2_s1_chipselect,                     --                                           .chipselect
			Hex_3_4_s1_address                               => mm_interconnect_0_hex_3_4_s1_address,                        --                                 Hex_3_4_s1.address
			Hex_3_4_s1_write                                 => mm_interconnect_0_hex_3_4_s1_write,                          --                                           .write
			Hex_3_4_s1_readdata                              => mm_interconnect_0_hex_3_4_s1_readdata,                       --                                           .readdata
			Hex_3_4_s1_writedata                             => mm_interconnect_0_hex_3_4_s1_writedata,                      --                                           .writedata
			Hex_3_4_s1_chipselect                            => mm_interconnect_0_hex_3_4_s1_chipselect,                     --                                           .chipselect
			Hex_5_6_s1_address                               => mm_interconnect_0_hex_5_6_s1_address,                        --                                 Hex_5_6_s1.address
			Hex_5_6_s1_write                                 => mm_interconnect_0_hex_5_6_s1_write,                          --                                           .write
			Hex_5_6_s1_readdata                              => mm_interconnect_0_hex_5_6_s1_readdata,                       --                                           .readdata
			Hex_5_6_s1_writedata                             => mm_interconnect_0_hex_5_6_s1_writedata,                      --                                           .writedata
			Hex_5_6_s1_chipselect                            => mm_interconnect_0_hex_5_6_s1_chipselect,                     --                                           .chipselect
			JTAG_UART_avalon_jtag_slave_address              => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,       --                JTAG_UART_avalon_jtag_slave.address
			JTAG_UART_avalon_jtag_slave_write                => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,         --                                           .write
			JTAG_UART_avalon_jtag_slave_read                 => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,          --                                           .read
			JTAG_UART_avalon_jtag_slave_readdata             => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,      --                                           .readdata
			JTAG_UART_avalon_jtag_slave_writedata            => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,     --                                           .writedata
			JTAG_UART_avalon_jtag_slave_waitrequest          => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,   --                                           .waitrequest
			JTAG_UART_avalon_jtag_slave_chipselect           => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,    --                                           .chipselect
			leds_s1_address                                  => mm_interconnect_0_leds_s1_address,                           --                                    leds_s1.address
			leds_s1_write                                    => mm_interconnect_0_leds_s1_write,                             --                                           .write
			leds_s1_readdata                                 => mm_interconnect_0_leds_s1_readdata,                          --                                           .readdata
			leds_s1_writedata                                => mm_interconnect_0_leds_s1_writedata,                         --                                           .writedata
			leds_s1_chipselect                               => mm_interconnect_0_leds_s1_chipselect,                        --                                           .chipselect
			MUTEX_s1_address                                 => mm_interconnect_0_mutex_s1_address,                          --                                   MUTEX_s1.address
			MUTEX_s1_write                                   => mm_interconnect_0_mutex_s1_write,                            --                                           .write
			MUTEX_s1_read                                    => mm_interconnect_0_mutex_s1_read,                             --                                           .read
			MUTEX_s1_readdata                                => mm_interconnect_0_mutex_s1_readdata,                         --                                           .readdata
			MUTEX_s1_writedata                               => mm_interconnect_0_mutex_s1_writedata,                        --                                           .writedata
			MUTEX_s1_chipselect                              => mm_interconnect_0_mutex_s1_chipselect,                       --                                           .chipselect
			Processor1_debug_mem_slave_address               => mm_interconnect_0_processor1_debug_mem_slave_address,        --                 Processor1_debug_mem_slave.address
			Processor1_debug_mem_slave_write                 => mm_interconnect_0_processor1_debug_mem_slave_write,          --                                           .write
			Processor1_debug_mem_slave_read                  => mm_interconnect_0_processor1_debug_mem_slave_read,           --                                           .read
			Processor1_debug_mem_slave_readdata              => mm_interconnect_0_processor1_debug_mem_slave_readdata,       --                                           .readdata
			Processor1_debug_mem_slave_writedata             => mm_interconnect_0_processor1_debug_mem_slave_writedata,      --                                           .writedata
			Processor1_debug_mem_slave_byteenable            => mm_interconnect_0_processor1_debug_mem_slave_byteenable,     --                                           .byteenable
			Processor1_debug_mem_slave_waitrequest           => mm_interconnect_0_processor1_debug_mem_slave_waitrequest,    --                                           .waitrequest
			Processor1_debug_mem_slave_debugaccess           => mm_interconnect_0_processor1_debug_mem_slave_debugaccess,    --                                           .debugaccess
			Processor2_debug_mem_slave_address               => mm_interconnect_0_processor2_debug_mem_slave_address,        --                 Processor2_debug_mem_slave.address
			Processor2_debug_mem_slave_write                 => mm_interconnect_0_processor2_debug_mem_slave_write,          --                                           .write
			Processor2_debug_mem_slave_read                  => mm_interconnect_0_processor2_debug_mem_slave_read,           --                                           .read
			Processor2_debug_mem_slave_readdata              => mm_interconnect_0_processor2_debug_mem_slave_readdata,       --                                           .readdata
			Processor2_debug_mem_slave_writedata             => mm_interconnect_0_processor2_debug_mem_slave_writedata,      --                                           .writedata
			Processor2_debug_mem_slave_byteenable            => mm_interconnect_0_processor2_debug_mem_slave_byteenable,     --                                           .byteenable
			Processor2_debug_mem_slave_waitrequest           => mm_interconnect_0_processor2_debug_mem_slave_waitrequest,    --                                           .waitrequest
			Processor2_debug_mem_slave_debugaccess           => mm_interconnect_0_processor2_debug_mem_slave_debugaccess,    --                                           .debugaccess
			pushbutton_s1_address                            => mm_interconnect_0_pushbutton_s1_address,                     --                              pushbutton_s1.address
			pushbutton_s1_write                              => mm_interconnect_0_pushbutton_s1_write,                       --                                           .write
			pushbutton_s1_readdata                           => mm_interconnect_0_pushbutton_s1_readdata,                    --                                           .readdata
			pushbutton_s1_writedata                          => mm_interconnect_0_pushbutton_s1_writedata,                   --                                           .writedata
			pushbutton_s1_chipselect                         => mm_interconnect_0_pushbutton_s1_chipselect,                  --                                           .chipselect
			RAM1_s1_address                                  => mm_interconnect_0_ram1_s1_address,                           --                                    RAM1_s1.address
			RAM1_s1_write                                    => mm_interconnect_0_ram1_s1_write,                             --                                           .write
			RAM1_s1_readdata                                 => mm_interconnect_0_ram1_s1_readdata,                          --                                           .readdata
			RAM1_s1_writedata                                => mm_interconnect_0_ram1_s1_writedata,                         --                                           .writedata
			RAM1_s1_byteenable                               => mm_interconnect_0_ram1_s1_byteenable,                        --                                           .byteenable
			RAM1_s1_chipselect                               => mm_interconnect_0_ram1_s1_chipselect,                        --                                           .chipselect
			RAM1_s1_clken                                    => mm_interconnect_0_ram1_s1_clken,                             --                                           .clken
			RAM2_s1_address                                  => mm_interconnect_0_ram2_s1_address,                           --                                    RAM2_s1.address
			RAM2_s1_write                                    => mm_interconnect_0_ram2_s1_write,                             --                                           .write
			RAM2_s1_readdata                                 => mm_interconnect_0_ram2_s1_readdata,                          --                                           .readdata
			RAM2_s1_writedata                                => mm_interconnect_0_ram2_s1_writedata,                         --                                           .writedata
			RAM2_s1_byteenable                               => mm_interconnect_0_ram2_s1_byteenable,                        --                                           .byteenable
			RAM2_s1_chipselect                               => mm_interconnect_0_ram2_s1_chipselect,                        --                                           .chipselect
			RAM2_s1_clken                                    => mm_interconnect_0_ram2_s1_clken,                             --                                           .clken
			rooms_manager_0_avalon_slave_0_write             => mm_interconnect_0_rooms_manager_0_avalon_slave_0_write,      --             rooms_manager_0_avalon_slave_0.write
			rooms_manager_0_avalon_slave_0_writedata         => mm_interconnect_0_rooms_manager_0_avalon_slave_0_writedata,  --                                           .writedata
			rooms_manager_0_avalon_slave_0_chipselect        => mm_interconnect_0_rooms_manager_0_avalon_slave_0_chipselect, --                                           .chipselect
			SHARED_MEMORY_s1_address                         => mm_interconnect_0_shared_memory_s1_address,                  --                           SHARED_MEMORY_s1.address
			SHARED_MEMORY_s1_write                           => mm_interconnect_0_shared_memory_s1_write,                    --                                           .write
			SHARED_MEMORY_s1_readdata                        => mm_interconnect_0_shared_memory_s1_readdata,                 --                                           .readdata
			SHARED_MEMORY_s1_writedata                       => mm_interconnect_0_shared_memory_s1_writedata,                --                                           .writedata
			SHARED_MEMORY_s1_byteenable                      => mm_interconnect_0_shared_memory_s1_byteenable,               --                                           .byteenable
			SHARED_MEMORY_s1_chipselect                      => mm_interconnect_0_shared_memory_s1_chipselect,               --                                           .chipselect
			SHARED_MEMORY_s1_clken                           => mm_interconnect_0_shared_memory_s1_clken,                    --                                           .clken
			sw_sliders_s1_address                            => mm_interconnect_0_sw_sliders_s1_address,                     --                              sw_sliders_s1.address
			sw_sliders_s1_write                              => mm_interconnect_0_sw_sliders_s1_write,                       --                                           .write
			sw_sliders_s1_readdata                           => mm_interconnect_0_sw_sliders_s1_readdata,                    --                                           .readdata
			sw_sliders_s1_writedata                          => mm_interconnect_0_sw_sliders_s1_writedata,                   --                                           .writedata
			sw_sliders_s1_chipselect                         => mm_interconnect_0_sw_sliders_s1_chipselect,                  --                                           .chipselect
			Timer1_s1_address                                => mm_interconnect_0_timer1_s1_address,                         --                                  Timer1_s1.address
			Timer1_s1_write                                  => mm_interconnect_0_timer1_s1_write,                           --                                           .write
			Timer1_s1_readdata                               => mm_interconnect_0_timer1_s1_readdata,                        --                                           .readdata
			Timer1_s1_writedata                              => mm_interconnect_0_timer1_s1_writedata,                       --                                           .writedata
			Timer1_s1_chipselect                             => mm_interconnect_0_timer1_s1_chipselect,                      --                                           .chipselect
			Timer2_s1_address                                => mm_interconnect_0_timer2_s1_address,                         --                                  Timer2_s1.address
			Timer2_s1_write                                  => mm_interconnect_0_timer2_s1_write,                           --                                           .write
			Timer2_s1_readdata                               => mm_interconnect_0_timer2_s1_readdata,                        --                                           .readdata
			Timer2_s1_writedata                              => mm_interconnect_0_timer2_s1_writedata,                       --                                           .writedata
			Timer2_s1_chipselect                             => mm_interconnect_0_timer2_s1_chipselect                       --                                           .chipselect
		);

	irq_mapper : component Lab7_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			sender_irq    => processor1_irq_irq              --    sender.irq
		);

	irq_mapper_001 : component Lab7_irq_mapper_001
		port map (
			clk           => clk_clk,                            --       clk.clk
			reset         => rst_controller_002_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_001_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver0_irq,           -- receiver2.irq
			receiver3_irq => irq_mapper_receiver2_irq,           -- receiver3.irq
			sender_irq    => processor2_irq_irq                  --    sender.irq
		);

	rst_controller : component lab7_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => processor1_debug_reset_request_reset, -- reset_in0.reset
			reset_in1      => processor1_debug_reset_request_reset, -- reset_in1.reset
			clk            => clk_clk,                              --       clk.clk
			reset_out      => rst_controller_reset_out_reset,       -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,   --          .reset_req
			reset_req_in0  => '0',                                  -- (terminated)
			reset_req_in1  => '0',                                  -- (terminated)
			reset_in2      => '0',                                  -- (terminated)
			reset_req_in2  => '0',                                  -- (terminated)
			reset_in3      => '0',                                  -- (terminated)
			reset_req_in3  => '0',                                  -- (terminated)
			reset_in4      => '0',                                  -- (terminated)
			reset_req_in4  => '0',                                  -- (terminated)
			reset_in5      => '0',                                  -- (terminated)
			reset_req_in5  => '0',                                  -- (terminated)
			reset_in6      => '0',                                  -- (terminated)
			reset_req_in6  => '0',                                  -- (terminated)
			reset_in7      => '0',                                  -- (terminated)
			reset_req_in7  => '0',                                  -- (terminated)
			reset_in8      => '0',                                  -- (terminated)
			reset_req_in8  => '0',                                  -- (terminated)
			reset_in9      => '0',                                  -- (terminated)
			reset_req_in9  => '0',                                  -- (terminated)
			reset_in10     => '0',                                  -- (terminated)
			reset_req_in10 => '0',                                  -- (terminated)
			reset_in11     => '0',                                  -- (terminated)
			reset_req_in11 => '0',                                  -- (terminated)
			reset_in12     => '0',                                  -- (terminated)
			reset_req_in12 => '0',                                  -- (terminated)
			reset_in13     => '0',                                  -- (terminated)
			reset_req_in13 => '0',                                  -- (terminated)
			reset_in14     => '0',                                  -- (terminated)
			reset_req_in14 => '0',                                  -- (terminated)
			reset_in15     => '0',                                  -- (terminated)
			reset_req_in15 => '0'                                   -- (terminated)
		);

	rst_controller_001 : component lab7_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 3,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => processor1_debug_reset_request_reset,   -- reset_in0.reset
			reset_in1      => processor2_debug_reset_request_reset,   -- reset_in1.reset
			reset_in2      => processor1_debug_reset_request_reset,   -- reset_in2.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_002 : component lab7_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => processor1_debug_reset_request_reset,   -- reset_in0.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_002_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_003 : component lab7_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => processor1_debug_reset_request_reset,   -- reset_in0.reset
			reset_in1      => processor2_debug_reset_request_reset,   -- reset_in1.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_003_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_sw_sliders_s1_write_ports_inv <= not mm_interconnect_0_sw_sliders_s1_write;

	mm_interconnect_0_timer1_s1_write_ports_inv <= not mm_interconnect_0_timer1_s1_write;

	mm_interconnect_0_pushbutton_s1_write_ports_inv <= not mm_interconnect_0_pushbutton_s1_write;

	mm_interconnect_0_timer2_s1_write_ports_inv <= not mm_interconnect_0_timer2_s1_write;

	mm_interconnect_0_hex_5_6_s1_write_ports_inv <= not mm_interconnect_0_hex_5_6_s1_write;

	mm_interconnect_0_hex_3_4_s1_write_ports_inv <= not mm_interconnect_0_hex_3_4_s1_write;

	mm_interconnect_0_hex_1_2_s1_write_ports_inv <= not mm_interconnect_0_hex_1_2_s1_write;

	mm_interconnect_0_leds_s1_write_ports_inv <= not mm_interconnect_0_leds_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

	rst_controller_003_reset_out_reset_ports_inv <= not rst_controller_003_reset_out_reset;

end architecture rtl; -- of Lab7
